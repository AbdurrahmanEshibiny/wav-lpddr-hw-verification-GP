// import wav_DFI_pkg::*;
`include "wddr_config.sv"
`include "wav_DFI_transfer.sv"

class wav_DFI_driver extends uvm_driver;
// use default value to adhere to the wavious standard, not #(wav_DFI_transfer); 

    wav_DFI_vif vif;
    uvm_phase driver_run_phase;
    wddr_config cfg;
	
    `uvm_component_utils_begin(wav_DFI_driver)
    `uvm_component_utils_end

    function new (string name = "wav_DFI_driver", uvm_component parent=null);
        super.new(name, parent);
        // FIXME: we need to solve the cfg problem
        uvm_config_db#(wddr_config)::get(null, "*", "cfg_obj", cfg);
    endfunction

    // function void connect_phase(uvm_phase phase);
        
    // endfunction

    virtual task run_phase(uvm_phase phase);
        driver_run_phase = phase;
        
        fork
            get_and_drive();
            respond_to_phyupd();
            respond_to_phymstr();
        join
    endtask
	
    virtual protected task get_and_drive();
        forever begin
            `uvm_info(get_type_name(), "wav_DFI driver waiting for the next item", UVM_MEDIUM);
            seq_item_port.get_next_item(req);
			`uvm_info(get_type_name(), "wav_DFI driver received the next item", UVM_MEDIUM);
			
            $cast(rsp, req.clone());

            rsp.set_id_info(req);
            `uvm_info(get_type_name(),$psprintf("wav_DFI driver start driving transfer :\n%s", rsp.sprint()), UVM_MEDIUM);

            drive_transaction(rsp);
            `uvm_info(get_type_name(),$psprintf("wav_DFI driver done driving transfer :\n%s", rsp.sprint()), UVM_MEDIUM);

			seq_item_port.item_done();
			seq_item_port.put_response(rsp);
        end
      endtask

    /*should we drive the signal through sequencer*/
      
    //reset tasks
    task automatic reset_lp(bit is_ctrl);
        if (is_ctrl) begin
            vif.mp_drv.cb_drv.lp_ctrl_req <= 0; 
            vif.mp_drv.cb_drv.lp_ctrl_wakeup <= 0; 
        end
        else begin
            vif.mp_drv.cb_drv.lp_data_req <= 0; 
            vif.mp_drv.cb_drv.lp_data_wakeup <= 0; 
        end
        `uvm_info(get_name(), "done resetting lp", UVM_MEDIUM);  
    endtask

    //drive lp interface according to the specified transaction
    task automatic drive_lp(wav_DFI_lp_transfer trans);  
        `uvm_info(get_name(), "Driving lp", UVM_MEDIUM);  
        @(posedge vif.mp_drv.cb_drv) 
        if (trans.is_ctrl) begin 
            vif.mp_drv.cb_drv.lp_ctrl_req <= trans.req; 
            vif.mp_drv.cb_drv.lp_ctrl_wakeup <= trans.wakeup; 
        end 
        else begin         
            vif.mp_drv.cb_drv.lp_data_req <= trans.req;         
            vif.mp_drv.cb_drv.lp_data_wakeup <= trans.wakeup; 
        end
        `uvm_info(get_name(), "done driving lp", UVM_MEDIUM);  

        if (trans.cyclesCount > 0) begin
            repeat (trans.cyclesCount) @(posedge vif.mp_drv.cb_drv);
            reset_lp(trans.is_ctrl);
        end
        `uvm_info(get_name(), "done driving lp transaction", UVM_MEDIUM);  
    endtask                        
        
    //drive ctrlupd interface according to the specified transaction
    task automatic drive_ctrlupd(wav_DFI_update_transfer trans);   
		int timer = 0;
        `uvm_info(get_name(), "Driving ctrlupd", UVM_MEDIUM);              
        @(posedge vif.mp_drv.cb_drv)         
        if (trans.is_ctrl) begin
            vif.mp_drv.cb_drv.ctrlupd_req <= trans.req;       
            `uvm_info(get_name(), "done driving ctrlupd", UVM_MEDIUM);  
            // if (trans.cyclesCount > 0) begin
            
			`uvm_info(get_name(), "wait for ctrlupd_ack goes HIGH", UVM_MEDIUM);
			forever begin
				@(posedge vif.mp_drv.cb_drv);
				++timer;
				if (vif.mp_drv.cb_drv.ctrlupd_ack == 1)
					break;
			end
            //wait(vif.mp_drv.cb_drv.ctrlupd_ack == 1);   
			`uvm_info(get_name(), "wait for ctrlupd_ack goes LOW, or timer to goes off", UVM_MEDIUM);
            //wait(vif.mp_drv.cb_drv.ctrlupd_ack == 0);
			forever begin
				@(posedge vif.mp_drv.cb_drv);
				++timer;
				if (vif.mp_drv.cb_drv.ctrlupd_ack == 0 || timer >= trans.cyclesCount)
					break;
			end
			
			vif.mp_drv.cb_drv.ctrlupd_req <= 0;
			`uvm_info(get_name(), "done resetting ctrlupd", UVM_MEDIUM);  
            // repeat(trans.cyclesCount) @(posedge vif.mp_drv.cb_drv);
            // vif.mp_drv.cb_drv.ctrlupd_req <= 0;
            // `uvm_info(get_name(), "Done resetting ctrlupd", UVM_MEDIUM); 
        end
    endtask

    task automatic drive_write(wav_DFI_write_transfer trans);  
        //trans.print();
        @(posedge vif.mp_drv.cb_drv);
            vif.mp_drv.cb_drv.dram_clk_disable[0] <= 0;
            vif.mp_drv.cb_drv.dram_clk_disable[1] <= 1;
            vif.mp_drv.cb_drv.dram_clk_disable[2] <= 1;
            vif.mp_drv.cb_drv.dram_clk_disable[3] <= 1;
            vif.mp_drv.cb_drv.cke[0] <= 2'b01;
            vif.mp_drv.cb_drv.cke[2] <= 2'b01;
            //wck
            vif.mp_drv.cb_drv.wck_cs[0] <= 2'b11; 
            vif.mp_drv.cb_drv.wck_cs[1] <= 2'b11;  
            vif.mp_drv.cb_drv.wck_cs[2] <= 2'b11; 
            vif.mp_drv.cb_drv.wck_cs[3] <= 2'b11;  
            vif.mp_drv.cb_drv.wck_en[0] <= 1; 
            vif.mp_drv.cb_drv.wck_en[1] <= 1;
            vif.mp_drv.cb_drv.wck_en[2] <= 1; 
            vif.mp_drv.cb_drv.wck_en[3] <= 1;
            vif.mp_drv.cb_drv.wck_toggle[0] <= 2'b01;
            vif.mp_drv.cb_drv.wck_toggle[1] <= 2'b01;
            vif.mp_drv.cb_drv.wck_toggle[2] <= 2'b01;
            vif.mp_drv.cb_drv.wck_toggle[3] <= 2'b01;
            
        @(posedge vif.mp_drv.cb_drv);
            //ACT1
            vif.mp_drv.cb_drv.address[0] <= 14'b0000000_0000111;
            vif.mp_drv.cb_drv.address[2] <= 14'b0000000_0000000;
            // cs
            vif.mp_drv.cb_drv.cs[0] <= 2'b01;
            vif.mp_drv.cb_drv.cs[2] <= 2'b01;
        @(posedge vif.mp_drv.cb_drv);
            //ACT2
            vif.mp_drv.cb_drv.address[0] <= 14'b0000000_0000011;
            vif.mp_drv.cb_drv.address[2] <= 14'b0000000_0000000;
        @(posedge vif.mp_drv.cb_drv);
            //CAS_WR
            vif.mp_drv.cb_drv.address[0] <= 14'b0000000_0011100;
            vif.mp_drv.cb_drv.address[2] <= 14'b0000000_0000000;
            
        @(posedge vif.mp_drv.cb_drv);
            //WR32
            vif.mp_drv.cb_drv.address[0] <= 14'b0000000_0000100;
            vif.mp_drv.cb_drv.address[2] <= 14'b0000000_1000000;
            //wck
            vif.mp_drv.cb_drv.wck_toggle[0] <= 2'b10;
            vif.mp_drv.cb_drv.wck_toggle[1] <= 2'b10;
            vif.mp_drv.cb_drv.wck_toggle[2] <= 2'b10;
            vif.mp_drv.cb_drv.wck_toggle[3] <= 2'b10;
        @(posedge vif.mp_drv.cb_drv);
            vif.mp_drv.cb_drv.wrdata_en[0] <= 1;
            vif.mp_drv.cb_drv.wrdata_en[1] <= 1;
            vif.mp_drv.cb_drv.wrdata_en[2] <= 1;
            vif.mp_drv.cb_drv.wrdata_en[3] <= 1;
            vif.mp_drv.cb_drv.wrdata[0] <= 64'habcd_ef98_1234_5678;
            vif.mp_drv.cb_drv.wrdata[2] <= 64'h1234_5678_abcd_ef98;
            vif.mp_drv.cb_drv.wrdata_cs[0] <= 2'b01;
            vif.mp_drv.cb_drv.wrdata_cs[2] <= 2'b01;
            
            
            
            vif.mp_drv.cb_drv.cs[0] <= 2'b00;
            vif.mp_drv.cb_drv.cs[2] <= 2'b00;
            vif.mp_drv.cb_drv.address[0] <= 14'b0000000_0000000;
            vif.mp_drv.cb_drv.address[2] <= 14'b0000000_0000000;


           #100ns;
           
        
           
        // @(posedge vif.mp_drv.cb_drv);
        //     //DES
        //     vif.mp_drv.cb_drv.address[0] <= 14'b0000000_0000000;
        
            
            //vif.mp_drv.cb_drv.parity_in[0] <= trans.parity_in[0]; 
               
            //vif.mp_drv.cb_drv.wrdata_mask[0] <= trans.wrdata_mask[0]; 
            
            //vif.mp_drv.cb_drv.dram_clk_disable[0] <= trans.dram_clk_disable[0];
            
            //vif.mp_drv.cb_drv.cke[0] <= trans.cke[0];
            
            
        // @(posedge vif.mp_drv.cb_drv);
        //     vif.mp_drv.cb_drv.address[0] <= 14'b0;
        //     vif.mp_drv.cb_drv.wrdata[0] <= 64'b0;
        //     //vif.mp_drv.cb_drv.parity_in[0] <= trans.parity_in[0]; 
        //     vif.mp_drv.cb_drv.wrdata_en[0] <= 0;   
        //     //vif.mp_drv.cb_drv.wrdata_mask[0] <= trans.wrdata_mask[0]; 
        //     vif.mp_drv.cb_drv.wck_cs[0] <= 2'b00;  
        //     vif.mp_drv.cb_drv.wck_en[0] <= 0; 
        //     vif.mp_drv.cb_drv.wck_toggle[0] <= 2'b00;
        //     vif.mp_drv.cb_drv.dram_clk_disable[0] <= 1;
        //     vif.mp_drv.cb_drv.wrdata_cs[0] <= 2'b00; 
        //     vif.mp_drv.cb_drv.cke[0] <= 0;
        //     vif.mp_drv.cb_drv.cs[0] <= 2'b00;
        
        
          
    endtask

    task automatic drive_status(wav_DFI_status_transfer trans);
        string msg;
        string freq_details;
        int tinit_start;
        vif.cb_drv.init_start <= 0;
        vif.cb_drv.freq_fsp <= trans.freq_fsp;
        vif.cb_drv.freq_ratio <= trans.freq_ratio;
        vif.cb_drv.frequency <= trans.frequency;
        @(vif.cb_drv);

        while (!vif.cb_drv.init_complete);
        vif.cb_drv.init_start <= 1;

        freq_details = $sformatf (
            "Frequency# = %0d, ", trans.frequency,
            "Freq Ratio = %0d, ", trans.freq_ratio,
            "FSP# = %0d", trans.freq_fsp
        );
        tinit_start = 1;

        while (tinit_start != 0) begin
            @(vif.cb_drv) begin
                if (vif.mp_drv.cb_drv.init_complete == 1'b0) begin
                    break;
                end
            end
            tinit_start++;
        end
        // vif.cb_drv.init_start <= 0;

        if (tinit_start == 0) begin
            msg = "PHY rejects new freq setting";
        end else begin
            msg = $sformatf (
                "PHY accepts new freq setting, tinit_start = %d", tinit_start);
        end
        `uvm_info (get_name(), {msg, "\n", freq_details}, UVM_MEDIUM)
        

        // need to drive dfi_cke and dfi_reset_n
        // until the dfi_init_complete signal is asserted.


        /*
        
        // FIXME: WE ARE TESTING FOR THE FREQUENCIES HERE
        // TODO: print the count of the timing if it succeeds
        */
    endtask

    // TODO: we need to declare variables for the current phase and the data
    // to be given to the signals on the command interface that are common
    // between read and write transactions (and any other transaction that
    // needs the command interface). These variables (could implemented as 
    // a struct) should be passed by reference as an input argument to the
    // drive_<sub_interface_name> task so that it can fill the struct
    // whenever the task needs to use the command interface. once the struct
    // is full (e.g., for a 4:1 system the struct contains 4 slices of command
    // interface signals) the task assigns the struct to the DFI interface. 
    // checking the fullness of the struct can be done by the current phase
    // variable.
    // Till now, the struct should consist of:
    // dfi_address, dfi_cke, dfi_cs,
    // dfi_dram_clk_disable, dfi_parity_in, dfi_reset

    // The above idea can be split into two main tasks:
    // task1: fills the command interface struct with the values it wants to
    // send
    // task2: whenever the struct has a size that is equal to or larger than
    // the frequency ratio. it assigns the values inside the struct to the
    // command interface. this can be used with other things as well

    // TODO: recheck that there are there are no other command interface
    // signals (other than the ones mentioned above) that are mentioned
    // in the DFI standard and implemented in the wavious design

    // TODO: we need to think about cases in ratioed systems when we want
    // to send multiple consecutive read instructions. the above idea
    // should solve it

    task drive_data (dfi_data_seq_item trans);
        // we will assume the frequency ratio is 1:1 for now
        // `uvm_info(get_name(), "Driving data", UVM_MEDIUM);
        data_trans curr_rw_item;
        data_trans next_rw_item;
        dfi_cmd_t cmd_;
        int rd_cmd_dly0;
        int rd_cmd_dly1;
        int j;
        for (j = 0; j < trans.data_items.size(); j++) begin
            curr_rw_item = trans.data_items[j];
            // write preamble to address bus
            foreach (curr_rw_item.preamble[i]) begin
                @(vif.mp_drv.cb_drv) begin
                    vif.mp_drv.cb_drv.address[0] <= curr_rw_item.preamble[i];
                end
            end
            // preamble done. choose which instruction to make
            if (curr_rw_item.dir == read_dir) begin
                cmd_ = DFI_RD16;
                cmd_[6:4] = curr_rw_item.address.col[5:3];
                cmd_[10:7] = curr_rw_item.address.ba;
                cmd_[12:11] = curr_rw_item.address.col[2:1];
                cmd_[3] = curr_rw_item.address.col[0];
                cmd_[13] = 1;
                if (j != (trans.data_items.size() - 1)) begin
                    next_rw_item = trans.data_items[j+1];
                end
                fork
                    begin
                        // write read instruction then NOP
                        // TODO: handle the problem of consectuive
                        // reads writes
                        @(vif.mp_drv.cb_drv) begin
                            vif.mp_drv.cb_drv.address[0] <= cmd_;                            
                        end
                        if (j == (trans.data_items.size() - 1)) begin
                            @(vif.mp_drv.cb_drv) begin
                                vif.mp_drv.cb_drv.address[0] <= DFI_NOP;
                            end
                        end else begin
                            if (next_rw_item.dir == read_dir) begin
                                rd_cmd_dly0 =
                                curr_rw_item.data_len
                                - next_rw_item.preamble.size() - 1;
                                if (rd_cmd_dly0 > 0) begin
                                    vif.mp_drv.cb_drv.address[0] <= DFI_NOP;
                                    repeat (rd_cmd_dly0) begin
                                        @(vif.mp_drv.cb_drv);
                                    end
                                end
                            end
                        end
                    end
                    begin
                        repeat (cfg.tphy_rdcslat) begin
                            @(vif.mp_drv.cb_drv);
                        end
                        vif.mp_drv.cb_drv.rddata_cs[0] <= curr_rw_item.cs;
                    end
                    begin
                        repeat (cfg.trddata_en) begin
                            @(vif.mp_drv.cb_drv);
                        end
                        vif.mp_drv.cb_drv.rddata_en[0] <= 1;
                        // cycles needed for rddata_en to stay 1
                        repeat (curr_rw_item.data_len) begin
                            @(vif.mp_drv.cb_drv);
                        end
                        if (j != (trans.data_items.size() - 1)) begin
                            next_rw_item = trans.data_items[j+1];
                            rd_cmd_dly1 =
                            curr_rw_item.data_len
                            - next_rw_item.preamble.size() - 1;
                            if (rd_cmd_dly1 < 0) begin
                                vif.mp_drv.cb_drv.rddata_en[0] <= 0;
                            end
                        end else begin
                            vif.mp_drv.cb_drv.rddata_en[0] <= 0;
                        end
                    end      
                join_any
            end
        end
    endtask

    //there are different types of DFI transactions 
    //this task checks the tr_type in the transaction and call the corresponding task 

    task automatic drive_transaction(wav_DFI_transfer trans);
        `uvm_info(get_name(), "write xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx", UVM_MEDIUM); 
        trans.print();
		fork begin
			wav_DFI_lp_transfer lp_trans;
			wav_DFI_update_transfer update_trans;
			wav_DFI_write_transfer write_trans;
            dfi_data_seq_item read_trans;
            wav_DFI_status_transfer status_trans;
		//add the remaining interface cases
			driver_run_phase.raise_objection(this, "start driving transaction");
			case(trans.tr_type)
				lp: begin
					$cast(lp_trans, trans);
					drive_lp(lp_trans);
				end 
				update: begin     
					$cast(update_trans, trans);
					drive_ctrlupd(update_trans); 
				end
				write: begin     
					$cast(write_trans, trans);
					drive_write(write_trans); 
				end
                status_freq: begin
                    $cast(status_trans, trans);
                    drive_status(status_trans);
                end
                data: begin
                    $cast(read_trans, trans);
                    drive_data(read_trans);
                end
			endcase
			driver_run_phase.drop_objection(this, "done driving transaction");
		end
        join_none
    endtask

    //monitors requests from the PHY on phyupd interface and grant them
    task automatic respond_to_phyupd();
        `uvm_info(get_name(), "starting respond_to_phyupd", UVM_MEDIUM);  
        forever begin
            @(posedge vif.mp_drv.cb_drv);
            if (vif.mp_drv.cb_drv.phyupd_req) begin
                driver_run_phase.raise_objection(this, "Respond to phyupd started");

                `uvm_info(get_name(), "Captured phyupd request HIGH", UVM_MEDIUM);  
                vif.mp_drv.cb_drv.phyupd_ack <= 1'b1;
                `uvm_info(get_name(), "Turned phyupd ack HIGH", UVM_MEDIUM);  

                wait(vif.mp_drv.cb_drv.phyupd_req == 0);

                `uvm_info(get_name(), "Captured phyupd request LOW", UVM_MEDIUM);  
                vif.mp_drv.cb_drv.phyupd_ack <= 1'b0;
                `uvm_info(get_name(), "Turned phyupd ack LOW", UVM_MEDIUM);  

                driver_run_phase.drop_objection(this, "Respond to phyupd finished");
            end
            else
                vif.mp_drv.cb_drv.phyupd_ack <= 1'b0;
        end
    endtask
    
    //monitors requests from the PHY on phymstr interface and grant them
    task automatic respond_to_phymstr();        
        `uvm_info(get_name(), "Waiting_to_phymstr", UVM_MEDIUM);   
        forever begin
            @(posedge vif.mp_drv.cb_drv) 
            if (vif.mp_drv.cb_drv.phymstr_req) begin 
                driver_run_phase.raise_objection(this, "Respond to phymstr started");

                `uvm_info(get_name(), "Captured phymstr request HIGH", UVM_MEDIUM);  
                vif.mp_drv.cb_drv.phymstr_ack <= 1'b1;
                `uvm_info(get_name(), "Turned phymstr ack HIGH", UVM_MEDIUM);
				
				wait(vif.mp_drv.cb_drv.phymstr_req == 0);
				
				`uvm_info(get_name(), "Captured phymstr request LOW", UVM_MEDIUM);  
                vif.mp_drv.cb_drv.phymstr_ack <= 1'b0;
                `uvm_info(get_name(), "Turned phymstr ack LOW", UVM_MEDIUM);

                driver_run_phase.drop_objection(this, "Respond to phymstr finished");
            end
            else
                vif.mp_drv.cb_drv.phymstr_ack <= 1'b0;
        end
    endtask

endclass