`include "DFI/DFI_agent/wav_DFI_transfer.sv"