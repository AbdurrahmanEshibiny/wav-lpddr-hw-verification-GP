`ifndef WAV_DFI_SEQ_LIB
`define WAV_DFI_SEQ_LIB

`include "uvm_macros.svh"
import uvm_pkg::*;

import wav_DFI_pkg::*;

`include "wav_DFI_ctrlupd_seq.sv"
`include "wav_DFI_lp_ctrl_seq.sv"
`include "wav_DFI_lp_data_seq.sv"

`endif