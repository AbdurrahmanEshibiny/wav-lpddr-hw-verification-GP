`include "DFI/DFI_agent/wav_DFI_transfer.sv"
`include "DFI/DFI_agent/wav_DFI_driver.sv"