`include "DFI/DFI_agent/wav_DFI_Agent_lib.svh"