typedef virtual wav_DFI_if wav_DFI_vif;