import uvm_pkg::*;

package wav_DFI_agent_pkg;

  `include "uvm_macros.svh"
  `include "DFI/DFI_agent/wav_DFI_defines.svh"
  `include "DFI/DFI_agent/wav_DFI_Agent_lib.svh"

endpackage