class wav_DFI_wck_seq extends uvm_sequence #(wav_DFI_wck_transfer);

    `uvm_object_utils(wav_DFI_wck_seq)

    function new(string name = "wav_DFI_wck_seq");
        super.new(name);  
    endfunction

   
endclass