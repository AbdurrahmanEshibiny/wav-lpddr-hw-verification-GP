`include "wav_DFI_ctrlupd_seq.sv"
`include "wav_DFI_lp_ctrl_seq.sv"
`include "wav_DFI_lp_data_seq.sv"