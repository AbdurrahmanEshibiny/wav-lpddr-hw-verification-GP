`include "DFI/DFI_agent/wav_DFI_Agent_lib.svh"
`include "DFI/sequences/wav_DFI_seq_lib.svh"