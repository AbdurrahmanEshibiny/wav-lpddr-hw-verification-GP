`ifndef WAV_DFI_SEQ_LIB
`define WAV_DFI_SEQ_LIB

`include "uvm_macros.svh"
import uvm_pkg::*;

import wav_DFI_pkg::*;


`endif