/*
TODO: the activation sequence (for read and write)
will be written here later on
*/