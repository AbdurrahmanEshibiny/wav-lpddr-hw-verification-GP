`ifndef WAV_DFI_SEQ_PKG_H_
`define WAV_DFI_SEQ_PKG_H_

package wav_DFI_SEQ_pkg;

  import uvm_pkg::*;

  import wav_DFI_pkg::*;

  `include "uvm_macros.svh"
  
  `include "DFI/sequences/wav_DFI_seq_lib.svh"

endpackage

`endif
