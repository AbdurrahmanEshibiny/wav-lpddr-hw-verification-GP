`include "DFI/DFI_agent/wav_DFI_if.sv"

package wav_DFI_pkg;
   import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "DFI/DFI_agent/wav_DFI_defines.svh"
  `include "DFI/wav_DFI_lib.svh"

endpackage