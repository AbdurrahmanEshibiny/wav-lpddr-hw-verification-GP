import uvm_pkg::*;

package wav_DFI_agent_pkg;

  `include "uvm_macros.svh"

endpackage